module servo_driver #(
    parameter integer FRAME_TICKS     = 1_000_000, // 20ms @ 50MHz
    parameter integer MIN_PULSE_TICK  = 50_000,    // 1.0ms @ 50MHz
    parameter integer MAX_PULSE_TICK  = 100_000,   // 2.0ms @ 50MHz
    // ���� ������ �̵��� ���� �Ķ���� �߰�
    parameter integer SLOW_TICK_MAX   = 5_000_000, // 0.1�� �ֱ�
    parameter integer STEP_SIZE_PULSE = 1000       // 0.1�ʸ��� �����̴� �޽� �� ũ�� (���� �ʿ�)
) (
    input  wire        clk,
    input  wire        rst,       
    input  wire [9:0]  duty_level,  // 0~1000. ���� ��ǥ ��Ƽ ���� (Target Duty)
    output wire        pwm_out
);
    
    // --- 1. ��������/���̾� ���� ---
    reg [19:0] cnt; // PWM ī���� (0~1,000,000-1)
    reg [22:0] slow_cnt; // 0.1�� Ÿ�̸�
    
    // ���� ���� �޽� ���� �����ϴ� �������� (���������� ��ǥ�� ������)
    reg [19:0] current_high_count; 
    
    // ��ǥ �޽� �� (���� ���� duty_level �Է¿� ��� ����)
    wire [19:0] target_high_count; 

    // --- 2. ��ǥ �޽� �� ��� (���� ��) ---
    // duty_level (0~1000)�� �޽� �� (50000~100000)���� ��ȯ
    assign target_high_count = MIN_PULSE_TICK +
                             ((MAX_PULSE_TICK - MIN_PULSE_TICK) * duty_level) / 1000;

    // --- 3. PWM ī���� (20ms ������) ---
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            cnt <= 20'd0;
        end else if (cnt == FRAME_TICKS - 1) begin
            cnt <= 20'd0;
        end else begin
            cnt <= cnt + 20'd1;
        end
    end

    // --- 4. ������ �̵� ���� (0.1�� �ֱ�) ---
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            slow_cnt <= 0;
            current_high_count <= MIN_PULSE_TICK; // �ʱ� ��ġ ����
        end else begin
            
            // 0.1�� Ÿ�̸� ������Ʈ
            if (slow_cnt == SLOW_TICK_MAX - 1) begin
                slow_cnt <= 0;
                
                // ��ǥ(target_high_count)�� ���� �޽� ��(current_high_count) ��
                if (current_high_count < target_high_count) begin
                    // ��ǥ���� ������ ���� (������ �̵�)
                    if (current_high_count + STEP_SIZE_PULSE > target_high_count)
                        current_high_count <= target_high_count; // ��ǥ �ʰ� ����
                    else
                        current_high_count <= current_high_count + STEP_SIZE_PULSE;
                        
                end else if (current_high_count > target_high_count) begin
                    // ��ǥ���� ũ�� ���� (���� �̵�)
                    if (current_high_count - STEP_SIZE_PULSE < target_high_count)
                        current_high_count <= target_high_count; // ��ǥ �ʰ� ����
                    else
                        current_high_count <= current_high_count - STEP_SIZE_PULSE;
                end
                
                // ��ǥ�� ������ ����
                
            end else begin
                slow_cnt <= slow_cnt + 1;
            end
        end
    end
    
    // --- 5. PWM ��� ---
    // ���� �޽� �� �������͸� ����Ͽ� PWM ��ȣ ����
    assign pwm_out = (cnt < current_high_count);

endmodule