module servo (
    input wire clk,       
    input wire rst,
    input wire l_ctrl,    
    input wire r_ctrl,    
    output wire servo     
);

parameter integer FRAME_TICK = 1000000; 
parameter integer PULSE_0   = 35000;   
parameter integer PULSE_180 = 115000; 
parameter integer STEP_SIZE = 2000;   


parameter integer SLOW_TICK_MAX = 5000000;

// �������� ����
reg [24:0] cnt;             // ������ ī���� (FRAME_TICK=1,000,000���� ī��Ʈ ����)
reg [24:0] target_pulse;    // ��ǥ �޽� �� �������� (PULSE_0 ~ PULSE_180 ���� ��)
reg [22:0] slow_cnt;        // �ӵ� ����� ī����

// --- target_pulse ���� ���� (�ӵ� ����) ---
always @(posedge clk or posedge rst) begin
    if (rst) begin
        slow_cnt <= 23'd0;
        target_pulse <= PULSE_0; 
    end
    else begin
        // 1. ���� Ŭ�� ī���� ������Ʈ
        if (slow_cnt == SLOW_TICK_MAX - 1) begin
            slow_cnt <= 23'd0; // ī���� ����
            
            // 2. 0.1�ʸ��� ��ư �Է� Ȯ�� �� target_pulse ������Ʈ
            if (r_ctrl) begin
                // ������ ��ư(r_ctrl) �޽��� ������ �� ����
                if (target_pulse + STEP_SIZE <= PULSE_180) begin
                    target_pulse <= target_pulse + STEP_SIZE;
                end else begin
                    target_pulse <= PULSE_180; // ���� ���� ����
                end
            end
            else if (l_ctrl) begin
                // ���� ��ư(l_ctrl) �޽��� ������ �� ����
                if (target_pulse - STEP_SIZE >= PULSE_0) begin
                    target_pulse <= target_pulse - STEP_SIZE;
                end else begin
                    target_pulse <= PULSE_0; // ���� ���� ����
                end
            end
        end
        else begin
            slow_cnt <= slow_cnt + 23'd1;
        end
    end
end

// --- PWM ������ �� ��� ���� ---
always @(posedge clk or posedge rst) begin
    if (rst) begin
        cnt <= 25'd0;
    end
    else begin
        if (cnt == FRAME_TICK - 1) begin // 20ms �ֱ� ����
            cnt <= 25'd0;
        end
        else begin
            cnt <= cnt + 25'd1;
        end
    end
end

// PWM ���: ī���Ͱ� ��ǥ �޽� ������ ���� �� High
assign servo = (cnt < target_pulse);

endmodule